library verilog;
use verilog.vl_types.all;
entity data_memory_tb is
end data_memory_tb;
