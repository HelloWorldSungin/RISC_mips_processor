module data_path_tb();
reg clk;
reg reset;
wire [31:0] writedata, dataadr;
wire memwrite;
// instantiate device to be tested
top dut (clk, reset, writedata, dataadr, memwrite);
// initialize test
initial
  begin
    reset <= 1; # 22; reset <= 0;
  end
// generate clock to sequence tests
always
  begin
    clk <=1; # 10; clk <= 0; # 10;
  end
// check results
/*
always @ (negedge clk)
  begin
    if (memwrite) begin
      if (dataadr === 29 & writedata === 19) begin
        $display ("Simulation succeeded");
        $stop;
      end else if (dataadr !== 28) begin
        $display ("Simulation failed");
        $stop;
      end
    end
  end
  */
endmodule
