
module ALU_control (input [1:0] ALUOp,
                    input [3:0] Opcode,
                    output reg [2:0] ALU_Cnt);

wire [5:0] ALUControl_In;
assign ALUControl_In = {ALUOp, Opcode};
always@(ALUControl_In)
  casex (ALUControl_In)
   6'b10xxxx: ALU_Cnt = 3'b000;
   6'b01xxxx: ALU_Cnt = 3'b001;
   6'b000010: ALU_Cnt = 3'b000;
   6'b000011: ALU_Cnt = 3'b001;
   6'b000100: ALU_Cnt = 3'b010;
   6'b000101: ALU_Cnt = 3'b011;
   6'b000110: ALU_Cnt = 3'b100;
   6'b000111: ALU_Cnt = 3'b101;
   6'b001000: ALU_Cnt = 3'b110;
   6'b001001: ALU_Cnt = 3'b111;
   default: ALU_Cnt = 3'b000;
  endcase
                       
 endmodule
