library verilog;
use verilog.vl_types.all;
entity inst_memory_tb is
end inst_memory_tb;
